`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/06/2025 10:06:44 AM
// Design Name: 
// Module Name: top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module top(
    
    input wclk,
    input rclk,
    input reset,
    input write_enable,
    input read_enable,
    input write_data_in,
    
    output fifo_occu_out,
    output fifo_occu_in,
    output full,
    output empty,
    output read_data_out
    );
    
    
    
    
    
    
    
    
    
    
endmodule



